module hamming_encoder (

    input logic [25 : 0] Din,

    output logic [31: 0] Dout

);



